module ddnf(
  input x1, x2, x3,
  output f1
);
  assign f1 = x1;
endmodule