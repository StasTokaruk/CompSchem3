library verilog;
use verilog.vl_types.all;
entity testbench_sum is
end testbench_sum;
