library verilog;
use verilog.vl_types.all;
entity tb_demux is
end tb_demux;
